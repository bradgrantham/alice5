
module Main(
    input wire clock,
    input wire reset_n,
    input wire run, // hold low and release reset to write inst and data
    output reg halted,

    input wire [15:0] ext_write_address,
    input wire [31:0] ext_write_data,
    input wire ext_enable_write_inst,
    input wire ext_enable_write_data,

    input wire ext_decode_inst,
    input wire [31:0] ext_inst_to_decode,
    output wire decode_opcode_is_branch,
    output wire decode_opcode_is_ALU_reg_imm,
    output wire decode_opcode_is_ALU_reg_reg,
    output wire decode_opcode_is_jal,
    output wire decode_opcode_is_jalr,
    output wire decode_opcode_is_lui,
    output wire decode_opcode_is_auipc,
    output wire decode_opcode_is_load,
    output wire decode_opcode_is_store,
    output wire decode_opcode_is_system,
    output wire decode_opcode_is_fadd,
    output wire decode_opcode_is_fsub,
    output wire decode_opcode_is_fmul,
    output wire decode_opcode_is_fdiv,
    output wire decode_opcode_is_fsgnj,
    output wire decode_opcode_is_fminmax,
    output wire decode_opcode_is_fsqrt,
    output wire decode_opcode_is_fcmp,
    output wire decode_opcode_is_fcvt_f2i,
    output wire decode_opcode_is_fmv_f2i,
    output wire decode_opcode_is_fcvt_i2f,
    output wire decode_opcode_is_fmv_i2f,
    output wire decode_opcode_is_flw,
    output wire decode_opcode_is_fsw,
    output wire decode_opcode_is_fmadd,
    output wire decode_opcode_is_fmsub,
    output wire decode_opcode_is_fnmsub,
    output wire decode_opcode_is_fnmadd,
    output wire [4:0] decode_rs1,
    output wire [4:0] decode_rs2,
    output wire [4:0] decode_rs3,
    output wire [4:0] decode_rd,
    output wire [1:0] decode_fmt,
    output wire [2:0] decode_funct3_rm,
    output wire [6:0] decode_funct7,
    output wire [4:0] decode_funct5,
    output wire [4:0] decode_shamt_ftype,
    output wire signed [11:0] decode_imm_alu_load,
    output wire signed [11:0] decode_imm_store,
    output wire signed [12:0] decode_imm_branch,
    output wire signed [31:0] decode_imm_upper,
    output wire signed [20:0] decode_imm_jump
);

    localparam WORD_WIDTH = 32;
    localparam REGISTER_ADDRESS_WIDTH = 5;
    localparam ADDRESS_WIDTH = 16;

    // CPU State Machine
    localparam STATE_INIT /* verilator public */ = 4'h00;
    localparam STATE_FETCH /* verilator public */ = 4'h01;
    localparam STATE_FETCH2 /* verilator public */ = 4'h02;
    localparam STATE_DECODE /* verilator public */ = 4'h03;
    localparam STATE_REGISTERS /* verilator public */ = 4'h04;
    localparam STATE_ALU /* verilator public */ = 4'h05;
    localparam STATE_STEPLOADSTORE /* verilator public */ = 4'h06;
    localparam STATE_HALTED /* verilator public */ = 4'h07;
    reg [3:0] state /* verilator public */;

    reg [WORD_WIDTH-1:0] PC /* verilator public */;

    // instruction latched for inst decoder
    reg [WORD_WIDTH-1:0] inst_to_decode /* verilator public */;

    // Instruction RAM write control
    reg [ADDRESS_WIDTH-1:0] inst_ram_address /* verilator public */;
    reg [WORD_WIDTH-1:0] inst_ram_in_data /* verilator public */;
    reg inst_ram_write;

    // Data RAM write control
    reg [ADDRESS_WIDTH-1:0] data_ram_address;
    reg [WORD_WIDTH-1:0] data_ram_in_data;
    reg data_ram_write;

    // Inst RAM read out
    wire [WORD_WIDTH-1:0] inst_ram_out_data /* verilator public */;

    // Data RAM read out
    wire [WORD_WIDTH-1:0] data_ram_out_data;

    BlockRam #(.WORD_WIDTH(32), .ADDRESS_WIDTH(ADDRESS_WIDTH))
        instRam(
            .clock(clock),
            .write_address({2'b00, inst_ram_address[ADDRESS_WIDTH-1:2]}),
            .write(inst_ram_write),
            .write_data(inst_ram_in_data),
            .read_address({2'b00, inst_ram_address[ADDRESS_WIDTH-1:2]}),
            .read_data(inst_ram_out_data));

    BlockRam #(.WORD_WIDTH(32), .ADDRESS_WIDTH(ADDRESS_WIDTH))
        dataRam(
            .clock(clock),
            .write_address({2'b00, data_ram_address[ADDRESS_WIDTH-1:2]}),
            .write(data_ram_write),
            .write_data(data_ram_in_data),
            .read_address({2'b00, data_ram_address[ADDRESS_WIDTH-1:2]}),
            .read_data(data_ram_out_data));

    wire [WORD_WIDTH-1:0] rs1_value /* verilator public */;
    wire [WORD_WIDTH-1:0] rs2_value /* verilator public */;
    reg [REGISTER_ADDRESS_WIDTH-1:0] rd_address;
    reg [WORD_WIDTH-1:0] alu_result;
    reg [WORD_WIDTH-1:0] rd_value;
    reg enable_write_rd;

    // Register bank.
    Registers registers(
        .clock(clock),

        .write_address(rd_address),
        .write(enable_write_rd),
        .write_data(rd_value),

        .read1_address(decode_rs1),
        .read1_data(rs1_value),

        .read2_address(decode_rs2),
        .read2_data(rs2_value));

    RISCVDecode #(.INSN_WIDTH(WORD_WIDTH))
        instDecode(
            .inst(inst_to_decode),
            .opcode_is_branch(decode_opcode_is_branch),
            .opcode_is_ALU_reg_imm(decode_opcode_is_ALU_reg_imm),
            .opcode_is_ALU_reg_reg(decode_opcode_is_ALU_reg_reg),
            .opcode_is_jal(decode_opcode_is_jal),
            .opcode_is_jalr(decode_opcode_is_jalr),
            .opcode_is_lui(decode_opcode_is_lui),
            .opcode_is_auipc(decode_opcode_is_auipc),
            .opcode_is_load(decode_opcode_is_load),
            .opcode_is_store(decode_opcode_is_store),
            .opcode_is_system(decode_opcode_is_system),
            .opcode_is_fadd(decode_opcode_is_fadd),
            .opcode_is_fsub(decode_opcode_is_fsub),
            .opcode_is_fmul(decode_opcode_is_fmul),
            .opcode_is_fdiv(decode_opcode_is_fdiv),
            .opcode_is_fsgnj(decode_opcode_is_fsgnj),
            .opcode_is_fminmax(decode_opcode_is_fminmax),
            .opcode_is_fsqrt(decode_opcode_is_fsqrt),
            .opcode_is_fcmp(decode_opcode_is_fcmp),
            .opcode_is_fcvt_f2i(decode_opcode_is_fcvt_f2i),
            .opcode_is_fmv_f2i(decode_opcode_is_fmv_f2i),
            .opcode_is_fcvt_i2f(decode_opcode_is_fcvt_i2f),
            .opcode_is_fmv_i2f(decode_opcode_is_fmv_i2f),
            .opcode_is_flw(decode_opcode_is_flw),
            .opcode_is_fsw(decode_opcode_is_fsw),
            .opcode_is_fmadd(decode_opcode_is_fmadd),
            .opcode_is_fmsub(decode_opcode_is_fmsub),
            .opcode_is_fnmsub(decode_opcode_is_fnmsub),
            .opcode_is_fnmadd(decode_opcode_is_fnmadd),
            .rs1(decode_rs1),
            .rs2(decode_rs2),
            .rs3(decode_rs3),
            .rd(decode_rd),
            .fmt(decode_fmt),
            .funct3_rm(decode_funct3_rm),
            .funct7(decode_funct7),
            .funct5(decode_funct5),
            .shamt_ftype(decode_shamt_ftype),
            .imm_alu_load(decode_imm_alu_load),
            .imm_store(decode_imm_store),
            .imm_branch(decode_imm_branch),
            .imm_upper(decode_imm_upper),
            .imm_jump(decode_imm_jump)
            );

    wire signed [WORD_WIDTH-1:0] alu_op1 /* verilator public */ ;
    wire signed [WORD_WIDTH-1:0] alu_op2 /* verilator public */ ;

    // If all parameters are signed, shorter parameters will be
    // sign-extended, according to Pong
    assign alu_op1 =
        (decode_opcode_is_ALU_reg_imm ||
           decode_opcode_is_ALU_reg_reg ||
           decode_opcode_is_jalr) ? $signed(rs1_value) :
        decode_opcode_is_lui ? $signed(decode_imm_upper) :
        decode_opcode_is_jal ? $signed(PC) :
        $signed(32'hdeadbeef);

    assign alu_op2 =
        (decode_opcode_is_ALU_reg_imm ||
            decode_opcode_is_jalr) ? decode_imm_alu_load :
        decode_opcode_is_ALU_reg_reg ? $signed(rs2_value) :
        decode_opcode_is_lui ? 0 :
        decode_opcode_is_jal ? $signed(decode_imm_jump) :
        $signed(32'hcafebabe);

    always @(posedge clock) begin
        if(!reset_n) begin

            state <= STATE_INIT;
            PC <= 0;
            inst_ram_write <= 0;
            data_ram_write <= 0;
            enable_write_rd <= 0;

            halted <= 0;

            // reset registers?  Could assume they're junk in the compiler and save gates

        end else begin

            if(!run) begin

                if(ext_decode_inst) begin
                    inst_to_decode <= ext_inst_to_decode;
                end

                if(ext_enable_write_inst) begin
                    inst_ram_address <= ext_write_address;
                    inst_ram_in_data <= ext_write_data;
                    inst_ram_write <= 1;
                end else begin
                    inst_ram_write <= 0;
                end

                if(ext_enable_write_data) begin
                    data_ram_address <= ext_write_address;
                    data_ram_in_data <= ext_write_data;
                    data_ram_write <= 1;
                end else begin
                    data_ram_write <= 0;
                end

            end else begin

                case (state)

                    STATE_INIT: begin
                        state <= STATE_FETCH;
                        PC <= 0;
                    end

                    STATE_FETCH: begin
                        // want PC to be settled here
                        // get instruction from memory[PC]
                        enable_write_rd <= 0;
                        inst_ram_address <= PC[15:0];
                        state <= STATE_FETCH2;
                        PC <= PC;
                    end

                    STATE_FETCH2: begin
                        state <= STATE_DECODE;
                    end

                    STATE_DECODE: begin
                        // clock the 32 bits of instruction into decoded signals
                        inst_to_decode <= inst_ram_out_data;
                        state <= STATE_REGISTERS;
                    end

                    STATE_REGISTERS: begin
                        halted <= decode_opcode_is_system &&
                            (decode_imm_alu_load[11:0] == 12'd1);
                        state <= STATE_ALU;
                    end

                    STATE_ALU: begin
                        // want decode of instruction and registers output to be settled here
                        // do ALU operation

                        // pretend all ops are add for now
                        alu_result <= alu_op1 + alu_op2;

                        rd_address <= decode_rd;

                        state <= halted ? STATE_HALTED : STATE_STEPLOADSTORE;
                    end

                    STATE_STEPLOADSTORE: begin
                        // want result of ALU to be settled here
                        // Would be output of ALU for branch and jalr or route from imm20 for branch

                        enable_write_rd <= (decode_opcode_is_ALU_reg_imm ||
                            decode_opcode_is_ALU_reg_reg ||
                            decode_opcode_is_lui ||
                            decode_opcode_is_jalr ||
                            decode_opcode_is_jal) &&
                            (rd_address != 0);
                        rd_value <= 
                            (decode_opcode_is_jalr || decode_opcode_is_jal) ? (PC + 4) :
                            $unsigned(alu_result);

			// We know the result of ALU for jal has
			// LSB 0, so just ignore LSB for both jal and
			// jalr
                        PC <= 
                            (decode_opcode_is_jal ||
                                 decode_opcode_is_jalr) ? $unsigned({alu_result[31:1],1'b0}) :
                            (PC + 4);

                        // load into registers?
                        // store from registers - need to stall reads from data, don't need to stall inst reads
                        state <= STATE_FETCH;
                    end

                    STATE_HALTED: begin
                        state <= STATE_HALTED;
                    end

                    default: begin
                        // error, just reset
                        state <= STATE_INIT;
                    end

                endcase
            end
        end
    end

endmodule
