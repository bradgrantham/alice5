
// Converts signed 32-bit int to 32-bit float.
module int_to_float(
    input wire [31:0] op,
    output wire [31:0] res);

// Make op positive.
wire sign = op[31];
wire [31:0] negative_op = -op;
wire [30:0] abs_op = op == 32'h80000000 ? 31'h7fffffff : sign ? negative_op[30:0] : op[30:0];

// Find the shift amount.
reg [4:0] shift;
always @(*) begin
    casex (abs_op)
        32'b1???????????????????????????????: shift = 5'd31;
        32'b01??????????????????????????????: shift = 5'd30;
        32'b001?????????????????????????????: shift = 5'd29;
        32'b0001????????????????????????????: shift = 5'd28;
        32'b00001???????????????????????????: shift = 5'd27;
        32'b000001??????????????????????????: shift = 5'd26;
        32'b0000001?????????????????????????: shift = 5'd25;
        32'b00000001????????????????????????: shift = 5'd24;
        32'b000000001???????????????????????: shift = 5'd23;
        32'b0000000001??????????????????????: shift = 5'd22;
        32'b00000000001?????????????????????: shift = 5'd21;
        32'b000000000001????????????????????: shift = 5'd20;
        32'b0000000000001???????????????????: shift = 5'd19;
        32'b00000000000001??????????????????: shift = 5'd18;
        32'b000000000000001?????????????????: shift = 5'd17;
        32'b0000000000000001????????????????: shift = 5'd16;
        32'b00000000000000001???????????????: shift = 5'd15;
        32'b000000000000000001??????????????: shift = 5'd14;
        32'b0000000000000000001?????????????: shift = 5'd13;
        32'b00000000000000000001????????????: shift = 5'd12;
        32'b000000000000000000001???????????: shift = 5'd11;
        32'b0000000000000000000001??????????: shift = 5'd10;
        32'b00000000000000000000001?????????: shift = 5'd9;
        32'b000000000000000000000001????????: shift = 5'd8;
        32'b0000000000000000000000001???????: shift = 5'd7;
        32'b00000000000000000000000001??????: shift = 5'd6;
        32'b000000000000000000000000001?????: shift = 5'd5;
        32'b0000000000000000000000000001????: shift = 5'd4;
        32'b00000000000000000000000000001???: shift = 5'd3;
        32'b000000000000000000000000000001??: shift = 5'd2;
        32'b0000000000000000000000000000001?: shift = 5'd1;
        32'b00000000000000000000000000000001: shift = 5'd0;
        32'b00000000000000000000000000000000: shift = 5'd0; // Doesn't matter, not used.
    endcase
end

wire is_zero = !|op;
wire [7:0] exp_part = 127 + shift;
wire [22:0] fract_part = shift < 23 ? abs_op << (23 - shift) : abs_op >> (shift - 23);
assign res = is_zero ? 32'h0 : { sign, exp_part, fract_part };

endmodule
